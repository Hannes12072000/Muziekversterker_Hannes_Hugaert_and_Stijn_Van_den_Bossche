Muziek versterker H&S
V1      57      0       DC      15
V2      58      0       DC      -15
V3      1       0       AC  	1
V4      9       0       AC  	1
V5		13		0		AC		1

R1      2       3       100k
R2      3       4       100k
R3      6       7       100k
R4      6       17      100k
R5      9       10      100k
R6      13      14      100k
R7      12      7       22k
R8      16      17      22k
R9      19      20      10k
R10     20      21      10k
R11     19      23      100k
R12     23      25      10k
R13     23      26      22k
R14     23      27      10k
R15     24      28      10k
R16     24      29      22k
R17     24      30      10k
R18     31      43      22k
R19     37      45      10k
R20     38      45      22k
R21     39      45      10k
R22     40      46      10k
R23     41      46      22k
R24     42      46      10k
R25     36      44      22k
R26     48      50      100*200
R27     47      49      100*200
R28     49      51      100
R29     50      54      100
R30     22      24      100k
.PARAM SET=.5
.STEP PARAM(SET) 0, 1,.2
X1  0  5  4   POT PARAMS: R=750 SET={SET}
X2  0  11 10  POT PARAMS: R=750 SET={SET}
X3  0  14 15  POT PARAMS: R=750 SET={SET}
X4  37 31 25  POT PARAMS: R=750 SET={SET}
X5  38 32 26  POT PARAMS: R=750 SET={SET}
X6  27 33 39  POT PARAMS: R=750 SET={SET}
X7  40 34 28  POT PARAMS: R=750 SET={SET}
X8  29 35 38  POT PARAMS: R=750 SET={SET}
X9  30 36 42  POT PARAMS: R=750 SET={SET}
X10 49 0  50  POT PARAMS: R=750 SET={SET}
X11 0  52 51  POT PARAMS: R=750 SET={SET}
X12 0  52 51  POT PARAMS: R=750 SET={SET}

*R41     5       0       RMOD 1

C1 	5 	6 	1�
C2 	11 	12 	1�
C3 	15 	16 	1�
C4 	25	37 	2.2�
C5 	26 	38 	2.2�
C6 	33 	43 	1.5n
C7 	32 	43 	6.8n
C8 	34 	44 	1.5n
C9  29 	41 	2.2�
C10 30 	42 	2.2�
C11 35 	44 	6.8n
C12 45 	47 	1�
C13 46 	48 	1�

C14 1 	2 	2.2�
C15 7 	8 	2.2�
C16 17 	18 	2.2�
C17 52 	55 	1�
C18 53 	56 	1�

X13  	0  		3  		57  	58  	4   	TL072
X14  	8  		19 		57  	58  	23  	TL072
X15  	18 		22 		57  	58  	24  	TL072
X16  	0  		43 		57  	58  	45   	TL072
X17  	0  		44 		57  	58  	46   	TL072


*//////////////////////////////////////////////////////////
*/ TL072 OPERATIONAL AMPLIFIER MACRO-MODEL
*//////////////////////////////////////////////////////////
* (REV N/A)      SUPPLY VOLTAGE: +/-15V
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OUTPUT
*                | | | | |
.SUBCKT TL072    1 2 3 4 5
*
  C1   11 12 3.498E-12
  C2    6  7 15.00E-12
  DC    5 53 DX
  DE   54  5 DX
  DLP  90 91 DX
  DLN  92 90 DX
  DP    4  3 DX
  EGND 99  0 POLY(2) (3,0) (4,0) 0 .5 .5
  FB    7 99 POLY(5) VB VC VE VLP VLN 0 4.715E6 -5E6 5E6 5E6 -5E6
  GA    6  0 11 12 282.8E-6
  GCM   0  6 10 99 8.942E-9
  ISS   3 10 DC 195.0E-6
  HLIM 90  0 VLIM 1K
  J1   11  2 10 JX
  J2   12  1 10 JX
  R2    6  9 100.0E3
  RD1   4 11 3.536E3
  RD2   4 12 3.536E3
  RO1   8  5 150
  RO2   7 99 150
  RP    3  4 2.143E3
  RSS  10 99 1.026E6
  VB    9  0 DC 0
  VC    3 53 DC 2.200
  VE   54  4 DC 2.200
  VLIM  7  8 DC 0
  VLP  91  0 DC 25
  VLN   0 92 DC 25
.MODEL DX D(IS=800.0E-18)
.MODEL JX PJF(IS=15.00E-12 BETA=270.1E-6 VTO=-1)
.ENDS

  	* This is the potentiometer
    *      _____
    *  1--|_____|--2
    *        |
    *        3
    
    *.SUBCKT potentiometer 1 2 3
    *.param w=limit(wiper,1m,.999)
    *R0 1 3 {R*(1-w)}
    *R1 3 2 {R*(w)}
    *.ENDS

.SUBCKT POT 1 T 2 PARAMS: VALUE=1K SET=0.5
RT 1 T {VALUE*(1-SET)+.001}
RB T 2 {VALUE*SET+.001}
.ENDS

*.model RMOD	RES(R=750)
*.STEP RES RMOD(R)	0, 750, 1500

.AC     dec     500     1       50k
.probe
.end